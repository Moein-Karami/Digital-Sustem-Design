module test #(parameter S) (input [S : 0]i, output [S : 0]o);
	assign o = i;
endmodule 